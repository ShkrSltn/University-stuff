LIBRARY ieee;
USE ieee.std_logic_1164.all; 
LIBRARY work;
ENTITY lab_2 IS 
	PORT
	(
		C :  IN  STD_LOGIC;
		Q0 :  OUT  STD_LOGIC;
		Q2 :  OUT  STD_LOGIC;
		Q1 :  OUT  STD_LOGIC;
		Q3 :  OUT  STD_LOGIC
	);
END lab_2;
ARCHITECTURE bdf_type OF lab_2 IS 
SIGNAL	SYNTHESIZED_WIRE_7 :  STD_LOGIC;
SIGNAL	DFF_inst :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_8 :  STD_LOGIC;
SIGNAL	DFF_inst2 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_9 :  STD_LOGIC;
SIGNAL	DFF_inst4 :  STD_LOGIC;
SIGNAL	SYNTHESIZED_WIRE_6 :  STD_LOGIC;
SIGNAL	DFF_inst6 :  STD_LOGIC;
BEGIN 
Q0 <= DFF_inst;
Q2 <= DFF_inst4;
Q1 <= DFF_inst2;
Q3 <= DFF_inst6;
PROCESS(C)
BEGIN
IF (RISING_EDGE(C)) THEN
	DFF_inst <= SYNTHESIZED_WIRE_7;
END IF;
END PROCESS;
SYNTHESIZED_WIRE_7 <= NOT(DFF_inst);
PROCESS(SYNTHESIZED_WIRE_7)
BEGIN
IF (RISING_EDGE(SYNTHESIZED_WIRE_7)) THEN
	DFF_inst2 <= SYNTHESIZED_WIRE_8;
END IF;
END PROCESS;
SYNTHESIZED_WIRE_8 <= NOT(DFF_inst2);
PROCESS(SYNTHESIZED_WIRE_8)
BEGIN
IF (RISING_EDGE(SYNTHESIZED_WIRE_8)) THEN
	DFF_inst4 <= SYNTHESIZED_WIRE_9;
END IF;
END PROCESS;
SYNTHESIZED_WIRE_9 <= NOT(DFF_inst4);
PROCESS(SYNTHESIZED_WIRE_9)
BEGIN
IF (RISING_EDGE(SYNTHESIZED_WIRE_9)) THEN
	DFF_inst6 <= SYNTHESIZED_WIRE_6;
END IF;
END PROCESS;
SYNTHESIZED_WIRE_6 <= NOT(DFF_inst6);
END bdf_type;
